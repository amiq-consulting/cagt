/******************************************************************************
 * (C) Copyright 2014 AMIQ Consulting
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * MODULE:      cagt_pkg.sv
 * PROJECT:     Common Agent
 * Description: This file contains all the includes of the cagt_pkg package.
 *******************************************************************************/

`ifndef CAGT_PKG_SV
	//protection against multiple includes
	`define CAGT_PKG_SV

	package cagt_pkg;
		import uvm_pkg::*;

		`include "uvm_macros.svh"

		`include "cagt_agent_config.sv"
		`include "cagt_coverage.sv"
		`include "cagt_monitor.sv"
		`include "cagt_driver.sv"
		`include "cagt_sequencer.sv"
		`include "cagt_agent.sv"

	endpackage

`endif
